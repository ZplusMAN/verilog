module demo ;
	function [7:0] getbyte ;
	endfunction 

	input [15:0] address ;
	begin 
	end
endmodule 
