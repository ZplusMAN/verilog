module demo;
	initial 
	begin 
		inputs = 'b000000;
		#10 inputs = b'011001;
		#10 inputs = b'000000;
	end
endmodule 
