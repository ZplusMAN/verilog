module demo;

	nand #10 nd1(a ,data, clock , clear );

endmodule 
