module demo;
	always @( posedge clock or posedge reset )
	begin 
	end 
endmodule 
