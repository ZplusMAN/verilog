module demo;
	task my_task ;
		input a , b ;
		inout c ;
		output d , e ;
		//执行任务相关的语句
		//

		c = foo1 ;
		d = foo2 ;
		e = foo3 ;
	endtask 
endmodule 

