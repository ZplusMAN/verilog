module demo;
	initial 
		$hello_verilog ;
endmodule 
