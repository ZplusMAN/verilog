module demo(input port1 , input port2 , output port3 , output  port4);

