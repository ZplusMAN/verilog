module top;
	initial 
	begin :block1 
		integer i ;
	end 
	initial 
	fork : block2 
		reg i ;
	join 

endmodule 
